`timescale 1ns/1ps

module scg_top (
  input 		 core_ddrc_core_clk,
  input 		 core_ddrc_rstn,


  output         io_As2ScgCmd_ready,
  input          io_As2ScgCmd_valid,
                 io_As2ScgCmd_bits_ADR_cmdtype,
                 io_As2ScgCmd_bits_ADR_adr_rank,
  input  [1:0]   io_As2ScgCmd_bits_ADR_adr_group,
                 io_As2ScgCmd_bits_ADR_adr_bank,
  input  [17:0]  io_As2ScgCmd_bits_ADR_adr_row,
  input  [9:0]   io_As2ScgCmd_bits_ADR_adr_col,
  input  [16:0]  io_As2ScgCmd_bits_ADR_adr_cmdToken,
  input          io_As2ScgCmd_bits_pri,
  input  [511:0] io_As2ScgWrdata_wdata,
  input  [63:0]  io_As2ScgWrdata_wstrb,
  input          io_Scg2AsRddata_ready,
  output         io_Scg2AsRddata_valid,
  output [511:0] io_Scg2AsRddata_bits_rdata,
  output [16:0]  io_Scg2AsRddata_bits_rtoken,
  input  [5:0]   io_scgregio_tRRDS,
                 io_scgregio_tRRDL,
  input  [7:0]   io_scgregio_tFAW,
  input  [5:0]   io_scgregio_tRCD,
                 io_scgregio_tRP,
  input  [7:0]   io_scgregio_tCCDS,
                 io_scgregio_tCCDL,
                 io_scgregio_tWTRS,
                 io_scgregio_tWTRL,
                 io_scgregio_tRTW,
                 io_scgregio_tWR,
                 io_scgregio_tRTP,
                 io_scgregio_tRAS,
                 io_scgregio_AL,
                 io_scgregio_WL,
                 io_scgregio_RL,
                 io_scgregio_BL,
  input  [15:0]  io_scgregio_tREFI,
  input  [31:0]  io_scgregio_tZQINTVL,
  input  [11:0]  io_scgregio_tRFC,
  input  [7:0]   io_scgregio_tZQCS,
                 io_scgregio_tphyWrlat,
                 io_scgregio_tphyWrcslat,
                 io_scgregio_tphyWrdata,
                 io_scgregio_trddataEn,
                 io_scgregio_tphyRdcslat,
                 io_scgregio_tphyRdlat,
                 io_scgregio_wrOdtDelay,
                 io_scgregio_wrOdtHold,
                 io_scgregio_rdOdtDelay,
                 io_scgregio_rdOdtHold,
  input          io_scgregio_dfiMode,
  input  [8:0]   io_scgregio_clspgTmInit,
  input  [1:0]   io_scgregio_prePolicy,
  output [2:0]   io_scgregio_RGState_0,
                 io_scgregio_RGState_1,
                 io_scgregio_RGState_2,
                 io_scgregio_RGState_3,
                 io_scgregio_refState,
  input          io_scgregio_dfiInitStart,
  output         io_scgregio_dfiInitComplete,
                 io_scgregio_ddrInitEnd,
  input  [20:0]  io_scgregio_dramRstn,
  input  [10:0]  io_scgregio_postCke,
  input  [23:0]  io_scgregio_preCke,
  input  [7:0]   io_scgregio_mrs2other,
  input  [3:0]   io_scgregio_mrs2mrs,
  input  [11:0]  io_scgregio_zqinit,
  input  [15:0]  io_scgregio_mrs1,
                 io_scgregio_mrs0,
                 io_scgregio_mrs3,
                 io_scgregio_mrs2,
                 io_scgregio_mrs5,
                 io_scgregio_mrs4,
                 io_scgregio_mrs6,
  input  [5:0]   io_scgregio_cmdGear,
  input  [7:0]   io_scgregio_syncGear,
                 io_scgregio_gearHold,
                 io_scgregio_gearSetup,
  input          io_scgregio_blkTGeardown,
                 io_scgregio_geardownMode,
                 io_calDone 
   
);

scg_wrapper u_scg_wrapper(
.core_ddrc_core_clk                     (core_ddrc_core_clk),
.core_ddrc_rstn                         (core_ddrc_rstn),


.io_As2ScgCmd_ready                     (io_As2ScgCmd_ready),
.io_As2ScgCmd_valid                     (io_As2ScgCmd_valid),
.io_As2ScgCmd_bits_ADR_cmdtype          (io_As2ScgCmd_bits_ADR_cmdtype),
.io_As2ScgCmd_bits_ADR_adr_rank         (io_As2ScgCmd_bits_ADR_adr_rank),
.io_As2ScgCmd_bits_ADR_adr_group        (io_As2ScgCmd_bits_ADR_adr_group),
.io_As2ScgCmd_bits_ADR_adr_bank         (io_As2ScgCmd_bits_ADR_adr_bank),
.io_As2ScgCmd_bits_ADR_adr_row          (io_As2ScgCmd_bits_ADR_adr_row),
.io_As2ScgCmd_bits_ADR_adr_col          (io_As2ScgCmd_bits_ADR_adr_col),
.io_As2ScgCmd_bits_ADR_adr_cmdToken     (io_As2ScgCmd_bits_ADR_adr_cmdToken),
.io_As2ScgCmd_bits_pri                  (io_As2ScgCmd_bits_pri),
.io_As2ScgWrdata_wdata                  (io_As2ScgWrdata_wdata),
.io_As2ScgWrdata_wstrb                  (io_As2ScgWrdata_wstrb),
.io_Scg2AsRddata_ready                  (io_Scg2AsRddata_ready),
.io_Scg2AsRddata_valid                  (io_Scg2AsRddata_valid),
.io_Scg2AsRddata_bits_rdata             (io_Scg2AsRddata_bits_rdata),
.io_Scg2AsRddata_bits_rtoken            (io_Scg2AsRddata_bits_rtoken),
.io_scgregio_tRRDS                      (io_scgregio_tRRDS),
.io_scgregio_tRRDL                      (io_scgregio_tRRDL),
.io_scgregio_tFAW                       (io_scgregio_tFAW),
.io_scgregio_tRCD                       (io_scgregio_tRCD),
.io_scgregio_tRP                        (io_scgregio_tRP),
.io_scgregio_tCCDS                      (io_scgregio_tCCDS),
.io_scgregio_tCCDL                      (io_scgregio_tCCDL),
.io_scgregio_tWTRS                      (io_scgregio_tWTRS),
.io_scgregio_tWTRL                      (io_scgregio_tWTRL),
.io_scgregio_tRTW                       (io_scgregio_tRTW),
.io_scgregio_tWR                        (io_scgregio_tWR),
.io_scgregio_tRTP                       (io_scgregio_tRTP),
.io_scgregio_tRAS                       (io_scgregio_tRAS),
.io_scgregio_AL                         (io_scgregio_AL),
.io_scgregio_WL                         (io_scgregio_WL),
.io_scgregio_RL                         (io_scgregio_RL),
.io_scgregio_BL                         (io_scgregio_BL),
.io_scgregio_tREFI                      (io_scgregio_tREFI),
.io_scgregio_tZQINTVL                   (io_scgregio_tZQINTVL),
.io_scgregio_tRFC                       (io_scgregio_tRFC),
.io_scgregio_tZQCS                      (io_scgregio_tZQCS),
.io_scgregio_tphyWrlat                  (io_scgregio_tphyWrlat),
.io_scgregio_tphyWrcslat                (io_scgregio_tphyWrcslat),
.io_scgregio_tphyWrdata                 (io_scgregio_tphyWrdata),
.io_scgregio_trddataEn                  (io_scgregio_trddataEn),
.io_scgregio_tphyRdcslat                (io_scgregio_tphyRdcslat),
.io_scgregio_tphyRdlat                  (io_scgregio_tphyRdlat),
.io_scgregio_wrOdtDelay                 (io_scgregio_wrOdtDelay),
.io_scgregio_wrOdtHold                  (io_scgregio_wrOdtHold),
.io_scgregio_rdOdtDelay                 (io_scgregio_rdOdtDelay),
.io_scgregio_rdOdtHold                  (io_scgregio_rdOdtHold),
.io_scgregio_dfiMode                    (io_scgregio_dfiMode),
.io_scgregio_clspgTmInit                (io_scgregio_clspgTmInit),
.io_scgregio_prePolicy                  (io_scgregio_prePolicy),
.io_scgregio_RGState_0                  (io_scgregio_RGState_0),
.io_scgregio_RGState_1                  (io_scgregio_RGState_1),
.io_scgregio_RGState_2                  (io_scgregio_RGState_2),
.io_scgregio_RGState_3                  (io_scgregio_RGState_3),
.io_scgregio_refState                   (io_scgregio_refState),
.io_scgregio_dfiInitStart               (io_scgregio_dfiInitStart),
.io_scgregio_dfiInitComplete            (io_scgregio_dfiInitComplete),
.io_scgregio_ddrInitEnd                 (io_scgregio_ddrInitEnd),
.io_scgregio_dramRstn                   (io_scgregio_dramRstn),
.io_scgregio_postCke                    (io_scgregio_postCke),
.io_scgregio_preCke                     (io_scgregio_preCke),
.io_scgregio_mrs2other                  (io_scgregio_mrs2other),
.io_scgregio_mrs2mrs                    (io_scgregio_mrs2mrs),
.io_scgregio_zqinit                     (io_scgregio_zqinit),
.io_scgregio_mrs1                       (io_scgregio_mrs1),
.io_scgregio_mrs0                       (io_scgregio_mrs0),
.io_scgregio_mrs3                       (io_scgregio_mrs3),
.io_scgregio_mrs2                       (io_scgregio_mrs2),
.io_scgregio_mrs5                       (io_scgregio_mrs5),
.io_scgregio_mrs4                       (io_scgregio_mrs4),
.io_scgregio_mrs6                       (io_scgregio_mrs6),
.io_scgregio_cmdGear                    (io_scgregio_cmdGear),
.io_scgregio_syncGear                   (io_scgregio_syncGear),
.io_scgregio_gearHold                   (io_scgregio_gearHold),
.io_scgregio_gearSetup                  (io_scgregio_gearSetup),
.io_scgregio_blkTGeardown               (io_scgregio_blkTGeardown),
.io_scgregio_geardownMode               (io_scgregio_geardownMode),
.io_calDone                             (io_calDone)
);


endmodule